----------------------------------------------------------------------------------
-- Company:			EBS INK-JET SYSTEMS POLAND 
-- Engineer: 		TOMASZ GRONOWICZ
-- 
-- Create Date:    07:01:33 10/17/2007 
-- Design Name: 	 Printer control logic
-- Module Name:    BREAK_VOL - Behavioral 
-- Project Name:	 EBS7100	
-- Target Devices: XC3S200-4PQ208
-- Tool versions:		ISE 8.2.03i	
-- Description: 		Breaking voltage and frequency generation
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments:
--		Breaking voltage wave and amplitude is generated by ADC
-- 		Voltage is set by SPI - MOSI singal is common for whole SPI's conected to XILINX
--		SCK is dedicated for this module (when bit SPI_SC(3) is set then SPI clk is
--		transferred to the ADC SPI clk.
--		The wave is generated by signals BR_CLR and BR_NLOAD, where BR_NLOAD sets the
--		voltage value and BR_CLR sets 0 on the ADC output. Both signals are controled by
--		DROP_CLK, so on the ADC output we get the square wave with DROP_CLK frequency and
--		voltage set by processor
--
-- Revision 0.02
-- During SPI transmission NLOAD and NCLR signals are hold high
-- Output signal is not generated
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BREAK_VOL is
    Port ( 
						BR_DROP_CLK : in   STD_LOGIC;
						BR_F16MHZ 	: in   STD_LOGIC;
						BR_SPI_CS 	: in   STD_LOGIC;
						BR_SPI_SCK 	: in   STD_LOGIC;
						
						BR_NCLR 		: out  STD_LOGIC;
						BR_NLOAD 		: out  STD_LOGIC;
						BR_SCLK 		: out  STD_LOGIC
					);
end BREAK_VOL;

architecture Behavioral of BREAK_VOL is

signal NLOAD 	: std_logic := '1';
signal NLOAD_CLR : std_logic := '1';

signal NCLR		: std_logic := '1';
signal NCLR_CLR : std_logic := '1';

begin

--Generate NLOAD signal ----------------------------------------
NLOAD_PROC:process(BR_DROP_CLK,NLOAD_CLR)
begin
	if (NLOAD_CLR = '1') then
		NLOAD <= '1';
	elsif (BR_DROP_CLK'event and BR_DROP_CLK ='1') then
		NLOAD <= '0';
	end if;

end process NLOAD_PROC;

--Generate NCLR signal -----------------------------------------
NCLR_PROC:process(BR_DROP_CLK,NCLR_CLR)
begin
	if (NCLR_CLR = '1') then
		NCLR <= '1';
	elsif (BR_DROP_CLK'event and BR_DROP_CLK ='0') then
		NCLR <= '0';
	end if;

end process NCLR_PROC;

--Clear signals-------------------------------------------------
SIG_CLR:process(BR_F16MHZ)
begin
	if (BR_F16MHZ'event and BR_F16MHZ ='1') then
		if (NLOAD='0') then
			NLOAD_CLR <= '1';
		else
			NLOAD_CLR <= '0';
		end if;
		
		if (NCLR='0') then
			NCLR_CLR <= '1';
		else
			NCLR_CLR <= '0';
		end if;
		
	end if;
end process SIG_CLR;

BR_NLOAD <= '1' when (BR_SPI_CS='0') else NLOAD;
BR_NCLR  <= '1' when (BR_SPI_CS='0') else NCLR;

-- Re-direct SPI clk
BR_SCLK <= BR_SPI_SCK when (BR_SPI_CS='0') else '0';

end Behavioral;

